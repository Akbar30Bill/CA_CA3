
`timescale 1ns/1ns

module DataPath();
  
end
